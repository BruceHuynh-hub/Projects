module Multiplier (input [15:0] a, b, output [15:0] multOut);

	assign multOut = a * b;

endmodule
