module Adder (input [15:0] a, input [7:0] b, output [15:0] addOut);

	assign addOut = a + b;

endmodule
