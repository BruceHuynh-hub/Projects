module Adder (input [15:0] a, b, output [15:0] addOut);

	assign addOut = a + b;

endmodule
